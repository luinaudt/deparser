process($muxSel )
  begin  
    case $muxSel is
      $cases
    end process;
