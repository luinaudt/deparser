-------------------------------------------------------------------------------
-- Title      : axiStream
-- Project    : 
-------------------------------------------------------------------------------
-- File       : axiStream.vhdl
-- Author     : luinaud thomas  <luinaud@localhost.localdomain>
-- Company    : 
-- Created    : 2020-01-16
-- Last update: 2020-01-16
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: A simple AXI stream interface
-------------------------------------------------------------------------------
-- Copyright (c) 2020 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author          Description
-- 2020-01-16  1.0      Thomas Luinaud	Created
-------------------------------------------------------------------------------

