process($muxSel )
  begin  
    case $muxSel is
      $cases
    end case;
end process;
    
