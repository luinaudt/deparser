-------------------------------------------------------------------------------
-- Title      : axi stream
-- Project    : 
-------------------------------------------------------------------------------
--! \file       : axiStream_fifo.vhdl
--! \author     : luinaud thomas  <luinaud@localhost.localdomain>
--! \brief      : axi stream fifo to validate axi slave and master interface
-------------------------------------------------------------------------------
-- Company    : 
-- Created    : 2020-01-16
-- Last update: 2020-01-23
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: FIFO : Slave --> Master
-------------------------------------------------------------------------------
-- Copyright (c) 2020 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2020-01-16  1.0      luinaud Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity AXI_stream is

  generic (
    reset_polarity : std_logic := '0';   --! reset polartity
    data_width     : natural   := 256;   --! width of the data bus in bits
    depth          : natural   := 512);  --! fifo depth 

  port (
    clk     : in  std_logic;            -- axi clk
    reset_n : in  std_logic;            -- asynchronous reset (active low)
    -- master interface
    ready_m : in  std_logic;            --! slave ready
    tlast_m : out std_logic;            --! TLAST
    valid_m : out std_logic;            --! indicate the transfer is valid
    data_m  : out std_logic_vector(data_width - 1 downto 0);  --! master data
    -- slave interface
    valid_s : in  std_logic;            --! master output is valid
    tlast_s : in  std_logic;            --! TLAST
    ready_s : out std_logic;            --! ready to receive
    data_s  : in  std_logic_vector(data_width - 1 downto 0)   --! slave data
    );
end entity;

architecture behavioral of AXI_stream is

  type ram_type is array (0 to depth - 1) of std_logic_vector(1 + data_width - 1 downto 0);
  signal fifo : ram_type;               --! memory to store elements

  signal tlast_i_in, tlast_i_out : std_logic;  --! tlast internal signals
  signal data_out                : std_logic_vector(data_width - 1 downto 0);  --! out of memory
  signal data_in                 : std_logic_vector(data_width - 1 downto 0);  --! input of memory
  signal head, head_next         : unsigned(8 downto 0);  --! head of fifo
  signal tail, tail_next         : unsigned(8 downto 0);  --! tail of fifo

  signal almost_empty : std_logic;      --! only one element to read
  signal almost_full  : std_logic;      --! only one place still available
  signal full, empty  : std_logic;      --! FIFO state
  signal ready_i      : std_logic;      --! the fifo is ready to receive value
  signal valid_i      : std_logic;      --! the fifo generates a valid output
begin  -- architecture behavioral
  ready_s    <= ready_i;
  valid_m    <= valid_i;
-- internal data signals :
--      IN signals must be synchronous
  data_in    <= data_s;
  tlast_i_in <= tlast_s;
--      OUT signals must be synchronous
  data_m     <= data_out;
  tlast_m    <= tlast_i_out;

  process (clk, reset_n)
  begin
    if reset_n = reset_polarity then
      full         <= '0';
      empty        <= '1';
      almost_full  <= '0';
      almost_empty <= '0';
    elsif rising_edge(clk) then
      almost_empty <= '0';
      almost_full <= '0';
      full  <= full;
      empty <= empty;
      if head_next = tail then          -- only one place free
        almost_full <= '1';
      end if;
      if tail_next = head then          -- only one element left
        almost_empty <= '1';
      end if;

      -- full and empty signal management
      if head /= tail then
        full  <= '0';
        empty <= '0';
      end if;

      if head = tail and almost_empty = '1' then
        empty <= '1';
      end if;

      if head = tail and almost_full = '1' then
        full <= '1';
      end if;
    end if;
  end process;

  process(head, head_next, tail, tail_next, empty, full, almost_full, almost_empty)
  begin
    head_next <= head + 1;
    tail_next <= tail + 1;
    valid_i   <= '1';
    ready_i   <= '1';

    if (head = tail and almost_empty = '1') or empty = '1' then
      valid_i <= '0';
    end if;

    if (head = tail and almost_full = '1') or full = '1' then
      ready_i <= '0';
    end if;

  end process;


  --! process to write and read from the fifo
  ram_proc : process(clk, reset_n)
  begin
    if reset_n = reset_polarity then
      tail        <= (others => '0');
      head        <= (others => '0');
      data_out    <= (others => '0');
      tlast_i_out <= '0';
    elsif rising_edge(clk) then
      if (ready_i and valid_s) = '1' then
        fifo(to_integer(head)) <= tlast_i_in & data_in;
        head                   <= head_next;
      end if;
      if (valid_i and ready_m) = '1' then
        tail        <= tail_next;
        data_out    <= fifo(to_integer(tail))(data_width - 1 downto 0);
        tlast_i_out <= fifo(to_integer(tail))(data_width);
      else
        data_out    <= (others => '0');
        tlast_i_out <= '0';
      end if;
    end if;
  end process;



end architecture behavioral;
